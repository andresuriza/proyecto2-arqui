module procesador(input logic clk,
						input logic	[7:0] q,
						output logic [18:0] address);

endmodule