`timescale 10ns/1ps

module and_tb();

    logic [15:0] a, b, c;

    and_ dut (
        .a(a),
        .b(b),
        .c(c)
    );

    initial begin
        a = 16'd3;  // 0000 0000 0000 0011
        b = 16'd3;  // 0000 0000 0000 0011
        #1ns;

        a = 16'd21; // 0000 0000 0001 0101
        b = 16'd9;  // 0000 0000 0000 1001
        #1ns;

        a = 16'd8;  // 0000 0000 0000 1000
        b = 16'd1;  // 0000 0000 0000 0001
        #1ns;

        a = 16'd0;  // 0000 0000 0000 0000
        b = 16'd0;  // 0000 0000 0000 0000
        #1ns;

        a = 16'd1;  // 0000 0000 0000 0001
        b = 16'd1;  // 0000 0000 0000 0001
        #1ns;

        $stop;
    end
endmodule
