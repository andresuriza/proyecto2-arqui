module shiftLeft(a, c);
    input [15:0] a;
    output [15:0] c;

    assign c = a << 1;
endmodule